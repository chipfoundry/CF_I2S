
/*
	Copyright 2024-2025 ChipFoundry, a DBA of Umbralogic Technologies LLC.

	Original Copyright 2024 Efabless Corp.
	Author: Efabless Corp. (ip_admin@efabless.com)

	Licensed under the Apache License, Version 2.0 (the "License");
	you may not use this file except in compliance with the License.
	You may obtain a copy of the License at

	    http://www.apache.org/licenses/LICENSE-2.0

	Unless required by applicable law or agreed to in writing, software
	distributed under the License is distributed on an "AS IS" BASIS,
	WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
	See the License for the specific language governing permissions and
	limitations under the License.

*/

`timescale			1ns/1ns

`default_nettype        none

`define     CLK(clk, period)        initial clk = 0; always #(period/2) clk = !clk;
`define     RSTn(rst, clk, duration)     initial rst = 1'bx; initial #5 rst = 1'b0; initial begin #duration; @(posedge clk) rst = 1'b1; end

`timescale  1ns/1ps

module CF_I2S_tb;
    localparam      AW = 4;
    localparam      DW = 32;
    reg             clk = 0;
    reg             rst_n;
    wire            sd, sdo;
    wire            ws;
    wire            sck;

    reg             fifo_rd = 1'b0;
    reg             fifo_clr = 1'b0;
    reg             fifo_en = 1'b1;
    
    reg [AW-1:0]    fifo_level_threshold = 5;

    wire            fifo_full;
    wire [AW-1:0]   fifo_level;
    wire            fifo_level_above;
    wire [31:0]     fifo_rdata;

    reg [5:0]       sample_size = 18;    
    reg [7:0]       sck_prescaler = (10/2)-1;

    reg [31:0]      avg_threshold = 32'h00_01_00_00;
    wire            avg_flag;

    reg [7:0]       clkdiv;

    localparam      FREQDIV = 10;

    CF_I2S #(.DW(DW), .AW(AW)) MUV (
        .clk(clk),
        .rst_n(rst_n),
        .sdi(sd),
        //.sdo(sdo),
        .ws(ws),
        .sck(sck),

        .fifo_en(fifo_en),
        .fifo_rd(fifo_rd),
        .fifo_clr(fifo_clr),
        .fifo_level_threshold(fifo_level_threshold),
        .fifo_full(fifo_full),
        .fifo_level(fifo_level),
        .fifo_level_above(fifo_level_above),
        .fifo_rdata(fifo_rdata),

        .sign_extend(1'b1),
        .left_justified(1'b1),
        .sample_size(sample_size),
        .sck_prescaler(sck_prescaler),
        .avg_threshold(avg_threshold),
        .avg_flag(avg_flag),
        .channels(2'b11),
        .en(1'b1)
    );

    i2s_mic vip (
        .sck(sck),
        .sdo(sd),
        .ws(ws)
    );

    `CLK(clk, 100)
    `RSTn(rst_n, clk, 1000)

    initial begin
        $dumpfile("CF_I2S_tb.vcd");
        $dumpvars;
        #1_500_000 $finish;
    end

    initial begin
        @(posedge fifo_level_above);
        repeat(5) begin
            @(posedge clk);
            fifo_rd <= 1'b1;
            @(posedge clk);
            fifo_rd <= 1'b0;
        end        
    end


endmodule


